module fast_serial_project():





endmodule
//EOF
