// picorv32_soc_avalon.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module picorv32_soc_avalon (
		input  wire       clk_clk,                     //              clk.clk
		output wire [7:0] led_gpio_cyc1000_led_signal, // led_gpio_cyc1000.led_signal
		input  wire       reset_reset_n                //            reset.reset_n
	);

	wire         picorv32_avalon_0_avm_m0_waitrequest;              // mm_interconnect_0:picorv32_avalon_0_avm_m0_waitrequest -> picorv32_avalon_0:avm_m0_waitrequest
	wire  [31:0] picorv32_avalon_0_avm_m0_readdata;                 // mm_interconnect_0:picorv32_avalon_0_avm_m0_readdata -> picorv32_avalon_0:avm_m0_readdata
	wire  [31:0] picorv32_avalon_0_avm_m0_address;                  // picorv32_avalon_0:avm_m0_address -> mm_interconnect_0:picorv32_avalon_0_avm_m0_address
	wire         picorv32_avalon_0_avm_m0_read;                     // picorv32_avalon_0:avm_m0_read -> mm_interconnect_0:picorv32_avalon_0_avm_m0_read
	wire   [3:0] picorv32_avalon_0_avm_m0_byteenable;               // picorv32_avalon_0:avm_m0_byteenable -> mm_interconnect_0:picorv32_avalon_0_avm_m0_byteenable
	wire         picorv32_avalon_0_avm_m0_readdatavalid;            // mm_interconnect_0:picorv32_avalon_0_avm_m0_readdatavalid -> picorv32_avalon_0:avm_m0_readdatavalid
	wire         picorv32_avalon_0_avm_m0_write;                    // picorv32_avalon_0:avm_m0_write -> mm_interconnect_0:picorv32_avalon_0_avm_m0_write
	wire  [31:0] picorv32_avalon_0_avm_m0_writedata;                // picorv32_avalon_0:avm_m0_writedata -> mm_interconnect_0:picorv32_avalon_0_avm_m0_writedata
	wire         mm_interconnect_0_led_gpio_0_avs_s0_chipselect;    // mm_interconnect_0:led_gpio_0_avs_s0_chipselect -> led_gpio_0:avs_s0_chipselect
	wire  [31:0] mm_interconnect_0_led_gpio_0_avs_s0_readdata;      // led_gpio_0:avs_s0_readdata -> mm_interconnect_0:led_gpio_0_avs_s0_readdata
	wire         mm_interconnect_0_led_gpio_0_avs_s0_waitrequest;   // led_gpio_0:avs_s0_waitrequest -> mm_interconnect_0:led_gpio_0_avs_s0_waitrequest
	wire   [1:0] mm_interconnect_0_led_gpio_0_avs_s0_address;       // mm_interconnect_0:led_gpio_0_avs_s0_address -> led_gpio_0:avs_s0_address
	wire         mm_interconnect_0_led_gpio_0_avs_s0_read;          // mm_interconnect_0:led_gpio_0_avs_s0_read -> led_gpio_0:avs_s0_read
	wire   [3:0] mm_interconnect_0_led_gpio_0_avs_s0_byteenable;    // mm_interconnect_0:led_gpio_0_avs_s0_byteenable -> led_gpio_0:avs_s0_byteenable
	wire         mm_interconnect_0_led_gpio_0_avs_s0_readdatavalid; // led_gpio_0:avs_s0_readdatavalid -> mm_interconnect_0:led_gpio_0_avs_s0_readdatavalid
	wire         mm_interconnect_0_led_gpio_0_avs_s0_write;         // mm_interconnect_0:led_gpio_0_avs_s0_write -> led_gpio_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_led_gpio_0_avs_s0_writedata;     // mm_interconnect_0:led_gpio_0_avs_s0_writedata -> led_gpio_0:avs_s0_writedata
	wire         mm_interconnect_0_fpga_ram_s1_chipselect;          // mm_interconnect_0:fpga_ram_s1_chipselect -> fpga_ram:chipselect
	wire  [31:0] mm_interconnect_0_fpga_ram_s1_readdata;            // fpga_ram:readdata -> mm_interconnect_0:fpga_ram_s1_readdata
	wire   [9:0] mm_interconnect_0_fpga_ram_s1_address;             // mm_interconnect_0:fpga_ram_s1_address -> fpga_ram:address
	wire   [3:0] mm_interconnect_0_fpga_ram_s1_byteenable;          // mm_interconnect_0:fpga_ram_s1_byteenable -> fpga_ram:byteenable
	wire         mm_interconnect_0_fpga_ram_s1_write;               // mm_interconnect_0:fpga_ram_s1_write -> fpga_ram:write
	wire  [31:0] mm_interconnect_0_fpga_ram_s1_writedata;           // mm_interconnect_0:fpga_ram_s1_writedata -> fpga_ram:writedata
	wire         mm_interconnect_0_fpga_ram_s1_clken;               // mm_interconnect_0:fpga_ram_s1_clken -> fpga_ram:clken
	wire         mm_interconnect_0_fpga_rom_s1_chipselect;          // mm_interconnect_0:fpga_rom_s1_chipselect -> fpga_rom:chipselect
	wire  [31:0] mm_interconnect_0_fpga_rom_s1_readdata;            // fpga_rom:readdata -> mm_interconnect_0:fpga_rom_s1_readdata
	wire         mm_interconnect_0_fpga_rom_s1_debugaccess;         // mm_interconnect_0:fpga_rom_s1_debugaccess -> fpga_rom:debugaccess
	wire   [9:0] mm_interconnect_0_fpga_rom_s1_address;             // mm_interconnect_0:fpga_rom_s1_address -> fpga_rom:address
	wire   [3:0] mm_interconnect_0_fpga_rom_s1_byteenable;          // mm_interconnect_0:fpga_rom_s1_byteenable -> fpga_rom:byteenable
	wire         mm_interconnect_0_fpga_rom_s1_write;               // mm_interconnect_0:fpga_rom_s1_write -> fpga_rom:write
	wire  [31:0] mm_interconnect_0_fpga_rom_s1_writedata;           // mm_interconnect_0:fpga_rom_s1_writedata -> fpga_rom:writedata
	wire         mm_interconnect_0_fpga_rom_s1_clken;               // mm_interconnect_0:fpga_rom_s1_clken -> fpga_rom:clken
	wire         mm_interconnect_0_mutex_0_s1_chipselect;           // mm_interconnect_0:mutex_0_s1_chipselect -> mutex_0:chipselect
	wire  [31:0] mm_interconnect_0_mutex_0_s1_readdata;             // mutex_0:data_to_cpu -> mm_interconnect_0:mutex_0_s1_readdata
	wire   [0:0] mm_interconnect_0_mutex_0_s1_address;              // mm_interconnect_0:mutex_0_s1_address -> mutex_0:address
	wire         mm_interconnect_0_mutex_0_s1_read;                 // mm_interconnect_0:mutex_0_s1_read -> mutex_0:read
	wire         mm_interconnect_0_mutex_0_s1_write;                // mm_interconnect_0:mutex_0_s1_write -> mutex_0:write
	wire  [31:0] mm_interconnect_0_mutex_0_s1_writedata;            // mm_interconnect_0:mutex_0_s1_writedata -> mutex_0:data_from_cpu
	wire  [31:0] picorv32_avalon_0_inr_irq0_irq;                    // irq_mapper:sender_irq -> picorv32_avalon_0:inr_irq0_irq
	wire         rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [fpga_ram:reset, fpga_rom:reset, irq_mapper:reset, led_gpio_0:reset_reset, mm_interconnect_0:picorv32_avalon_0_reset_reset_bridge_in_reset_reset, mutex_0:reset_n, picorv32_avalon_0:reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                // rst_controller:reset_req -> [fpga_ram:reset_req, fpga_rom:reset_req, rst_translator:reset_req_in]

	picorv32_soc_avalon_fpga_ram fpga_ram (
		.clk        (clk_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_fpga_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_fpga_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_fpga_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_fpga_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_fpga_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_fpga_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_fpga_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	picorv32_soc_avalon_fpga_rom fpga_rom (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (mm_interconnect_0_fpga_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_fpga_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_fpga_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_fpga_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_fpga_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_fpga_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_fpga_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_fpga_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	led_gpio led_gpio_0 (
		.avs_s0_address       (mm_interconnect_0_led_gpio_0_avs_s0_address),       //   avs_s0.address
		.avs_s0_read          (mm_interconnect_0_led_gpio_0_avs_s0_read),          //         .read
		.avs_s0_readdata      (mm_interconnect_0_led_gpio_0_avs_s0_readdata),      //         .readdata
		.avs_s0_readdatavalid (mm_interconnect_0_led_gpio_0_avs_s0_readdatavalid), //         .readdatavalid
		.avs_s0_write         (mm_interconnect_0_led_gpio_0_avs_s0_write),         //         .write
		.avs_s0_writedata     (mm_interconnect_0_led_gpio_0_avs_s0_writedata),     //         .writedata
		.avs_s0_waitrequest   (mm_interconnect_0_led_gpio_0_avs_s0_waitrequest),   //         .waitrequest
		.avs_s0_byteenable    (mm_interconnect_0_led_gpio_0_avs_s0_byteenable),    //         .byteenable
		.avs_s0_chipselect    (mm_interconnect_0_led_gpio_0_avs_s0_chipselect),    //         .chipselect
		.clock_clk            (clk_clk),                                           //    clock.clk
		.reset_reset          (rst_controller_reset_out_reset),                    //    reset.reset
		.led                  (led_gpio_cyc1000_led_signal)                        // led_gpio.led_signal
	);

	picorv32_soc_avalon_mutex_0 mutex_0 (
		.reset_n       (~rst_controller_reset_out_reset),         // reset.reset_n
		.clk           (clk_clk),                                 //   clk.clk
		.chipselect    (mm_interconnect_0_mutex_0_s1_chipselect), //    s1.chipselect
		.data_from_cpu (mm_interconnect_0_mutex_0_s1_writedata),  //      .writedata
		.read          (mm_interconnect_0_mutex_0_s1_read),       //      .read
		.write         (mm_interconnect_0_mutex_0_s1_write),      //      .write
		.data_to_cpu   (mm_interconnect_0_mutex_0_s1_readdata),   //      .readdata
		.address       (mm_interconnect_0_mutex_0_s1_address)     //      .address
	);

	picorv32_avalon picorv32_avalon_0 (
		.avm_m0_address       (picorv32_avalon_0_avm_m0_address),       //   avm_m0.address
		.avm_m0_read          (picorv32_avalon_0_avm_m0_read),          //         .read
		.avm_m0_waitrequest   (picorv32_avalon_0_avm_m0_waitrequest),   //         .waitrequest
		.avm_m0_readdata      (picorv32_avalon_0_avm_m0_readdata),      //         .readdata
		.avm_m0_readdatavalid (picorv32_avalon_0_avm_m0_readdatavalid), //         .readdatavalid
		.avm_m0_write         (picorv32_avalon_0_avm_m0_write),         //         .write
		.avm_m0_writedata     (picorv32_avalon_0_avm_m0_writedata),     //         .writedata
		.avm_m0_byteenable    (picorv32_avalon_0_avm_m0_byteenable),    //         .byteenable
		.clock_clk            (clk_clk),                                //    clock.clk
		.reset_reset          (rst_controller_reset_out_reset),         //    reset.reset
		.inr_irq0_irq         (picorv32_avalon_0_inr_irq0_irq)          // inr_irq0.irq
	);

	picorv32_soc_avalon_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                           //                                     clk_0_clk.clk
		.picorv32_avalon_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // picorv32_avalon_0_reset_reset_bridge_in_reset.reset
		.picorv32_avalon_0_avm_m0_address                    (picorv32_avalon_0_avm_m0_address),                  //                      picorv32_avalon_0_avm_m0.address
		.picorv32_avalon_0_avm_m0_waitrequest                (picorv32_avalon_0_avm_m0_waitrequest),              //                                              .waitrequest
		.picorv32_avalon_0_avm_m0_byteenable                 (picorv32_avalon_0_avm_m0_byteenable),               //                                              .byteenable
		.picorv32_avalon_0_avm_m0_read                       (picorv32_avalon_0_avm_m0_read),                     //                                              .read
		.picorv32_avalon_0_avm_m0_readdata                   (picorv32_avalon_0_avm_m0_readdata),                 //                                              .readdata
		.picorv32_avalon_0_avm_m0_readdatavalid              (picorv32_avalon_0_avm_m0_readdatavalid),            //                                              .readdatavalid
		.picorv32_avalon_0_avm_m0_write                      (picorv32_avalon_0_avm_m0_write),                    //                                              .write
		.picorv32_avalon_0_avm_m0_writedata                  (picorv32_avalon_0_avm_m0_writedata),                //                                              .writedata
		.fpga_ram_s1_address                                 (mm_interconnect_0_fpga_ram_s1_address),             //                                   fpga_ram_s1.address
		.fpga_ram_s1_write                                   (mm_interconnect_0_fpga_ram_s1_write),               //                                              .write
		.fpga_ram_s1_readdata                                (mm_interconnect_0_fpga_ram_s1_readdata),            //                                              .readdata
		.fpga_ram_s1_writedata                               (mm_interconnect_0_fpga_ram_s1_writedata),           //                                              .writedata
		.fpga_ram_s1_byteenable                              (mm_interconnect_0_fpga_ram_s1_byteenable),          //                                              .byteenable
		.fpga_ram_s1_chipselect                              (mm_interconnect_0_fpga_ram_s1_chipselect),          //                                              .chipselect
		.fpga_ram_s1_clken                                   (mm_interconnect_0_fpga_ram_s1_clken),               //                                              .clken
		.fpga_rom_s1_address                                 (mm_interconnect_0_fpga_rom_s1_address),             //                                   fpga_rom_s1.address
		.fpga_rom_s1_write                                   (mm_interconnect_0_fpga_rom_s1_write),               //                                              .write
		.fpga_rom_s1_readdata                                (mm_interconnect_0_fpga_rom_s1_readdata),            //                                              .readdata
		.fpga_rom_s1_writedata                               (mm_interconnect_0_fpga_rom_s1_writedata),           //                                              .writedata
		.fpga_rom_s1_byteenable                              (mm_interconnect_0_fpga_rom_s1_byteenable),          //                                              .byteenable
		.fpga_rom_s1_chipselect                              (mm_interconnect_0_fpga_rom_s1_chipselect),          //                                              .chipselect
		.fpga_rom_s1_clken                                   (mm_interconnect_0_fpga_rom_s1_clken),               //                                              .clken
		.fpga_rom_s1_debugaccess                             (mm_interconnect_0_fpga_rom_s1_debugaccess),         //                                              .debugaccess
		.led_gpio_0_avs_s0_address                           (mm_interconnect_0_led_gpio_0_avs_s0_address),       //                             led_gpio_0_avs_s0.address
		.led_gpio_0_avs_s0_write                             (mm_interconnect_0_led_gpio_0_avs_s0_write),         //                                              .write
		.led_gpio_0_avs_s0_read                              (mm_interconnect_0_led_gpio_0_avs_s0_read),          //                                              .read
		.led_gpio_0_avs_s0_readdata                          (mm_interconnect_0_led_gpio_0_avs_s0_readdata),      //                                              .readdata
		.led_gpio_0_avs_s0_writedata                         (mm_interconnect_0_led_gpio_0_avs_s0_writedata),     //                                              .writedata
		.led_gpio_0_avs_s0_byteenable                        (mm_interconnect_0_led_gpio_0_avs_s0_byteenable),    //                                              .byteenable
		.led_gpio_0_avs_s0_readdatavalid                     (mm_interconnect_0_led_gpio_0_avs_s0_readdatavalid), //                                              .readdatavalid
		.led_gpio_0_avs_s0_waitrequest                       (mm_interconnect_0_led_gpio_0_avs_s0_waitrequest),   //                                              .waitrequest
		.led_gpio_0_avs_s0_chipselect                        (mm_interconnect_0_led_gpio_0_avs_s0_chipselect),    //                                              .chipselect
		.mutex_0_s1_address                                  (mm_interconnect_0_mutex_0_s1_address),              //                                    mutex_0_s1.address
		.mutex_0_s1_write                                    (mm_interconnect_0_mutex_0_s1_write),                //                                              .write
		.mutex_0_s1_read                                     (mm_interconnect_0_mutex_0_s1_read),                 //                                              .read
		.mutex_0_s1_readdata                                 (mm_interconnect_0_mutex_0_s1_readdata),             //                                              .readdata
		.mutex_0_s1_writedata                                (mm_interconnect_0_mutex_0_s1_writedata),            //                                              .writedata
		.mutex_0_s1_chipselect                               (mm_interconnect_0_mutex_0_s1_chipselect)            //                                              .chipselect
	);

	picorv32_soc_avalon_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (picorv32_avalon_0_inr_irq0_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
