// led_example.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module led_example (
		output wire       blinkt_led_serial_serial_clk,            //                 blinkt_led_serial.serial_clk
		output wire       blinkt_led_serial_serial_data,           //                                  .serial_data
		output wire       bytes_to_packets_in_bytes_stream_ready,  //  bytes_to_packets_in_bytes_stream.ready
		input  wire       bytes_to_packets_in_bytes_stream_valid,  //                                  .valid
		input  wire [7:0] bytes_to_packets_in_bytes_stream_data,   //                                  .data
		input  wire       clk_clk,                                 //                               clk.clk
		input  wire       packets_to_bytes_out_bytes_stream_ready, // packets_to_bytes_out_bytes_stream.ready
		output wire       packets_to_bytes_out_bytes_stream_valid, //                                  .valid
		output wire [7:0] packets_to_bytes_out_bytes_stream_data,  //                                  .data
		input  wire       reset_reset_n,                           //                             reset.reset_n
		output wire [7:0] simple_leds_leds                         //                       simple_leds.leds
	);

	wire  [31:0] master_avalon_master_readdata;                     // mm_interconnect_0:master_avalon_master_readdata -> master:readdata
	wire         master_avalon_master_waitrequest;                  // mm_interconnect_0:master_avalon_master_waitrequest -> master:waitrequest
	wire  [31:0] master_avalon_master_address;                      // master:address -> mm_interconnect_0:master_avalon_master_address
	wire         master_avalon_master_read;                         // master:read -> mm_interconnect_0:master_avalon_master_read
	wire   [3:0] master_avalon_master_byteenable;                   // master:byteenable -> mm_interconnect_0:master_avalon_master_byteenable
	wire         master_avalon_master_readdatavalid;                // mm_interconnect_0:master_avalon_master_readdatavalid -> master:readdatavalid
	wire         master_avalon_master_write;                        // master:write -> mm_interconnect_0:master_avalon_master_write
	wire  [31:0] master_avalon_master_writedata;                    // master:writedata -> mm_interconnect_0:master_avalon_master_writedata
	wire         mm_interconnect_0_simple_led_0_avs_s0_chipselect;  // mm_interconnect_0:simple_led_0_avs_s0_chipselect -> simple_led_0:avs_s0_chipselect
	wire  [31:0] mm_interconnect_0_simple_led_0_avs_s0_readdata;    // simple_led_0:avs_s0_readdata -> mm_interconnect_0:simple_led_0_avs_s0_readdata
	wire         mm_interconnect_0_simple_led_0_avs_s0_waitrequest; // simple_led_0:avs_s0_waitrequest -> mm_interconnect_0:simple_led_0_avs_s0_waitrequest
	wire   [3:0] mm_interconnect_0_simple_led_0_avs_s0_address;     // mm_interconnect_0:simple_led_0_avs_s0_address -> simple_led_0:avs_s0_address
	wire         mm_interconnect_0_simple_led_0_avs_s0_read;        // mm_interconnect_0:simple_led_0_avs_s0_read -> simple_led_0:avs_s0_read
	wire         mm_interconnect_0_simple_led_0_avs_s0_write;       // mm_interconnect_0:simple_led_0_avs_s0_write -> simple_led_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_simple_led_0_avs_s0_writedata;   // mm_interconnect_0:simple_led_0_avs_s0_writedata -> simple_led_0:avs_s0_writedata
	wire         mm_interconnect_0_blinkt_led_0_avs_s0_chipselect;  // mm_interconnect_0:blinkt_led_0_avs_s0_chipselect -> blinkt_led_0:avs_s0_chipselect
	wire  [31:0] mm_interconnect_0_blinkt_led_0_avs_s0_readdata;    // blinkt_led_0:avs_s0_readdata -> mm_interconnect_0:blinkt_led_0_avs_s0_readdata
	wire         mm_interconnect_0_blinkt_led_0_avs_s0_waitrequest; // blinkt_led_0:avs_s0_waitrequest -> mm_interconnect_0:blinkt_led_0_avs_s0_waitrequest
	wire   [3:0] mm_interconnect_0_blinkt_led_0_avs_s0_address;     // mm_interconnect_0:blinkt_led_0_avs_s0_address -> blinkt_led_0:avs_s0_address
	wire         mm_interconnect_0_blinkt_led_0_avs_s0_read;        // mm_interconnect_0:blinkt_led_0_avs_s0_read -> blinkt_led_0:avs_s0_read
	wire         mm_interconnect_0_blinkt_led_0_avs_s0_write;       // mm_interconnect_0:blinkt_led_0_avs_s0_write -> blinkt_led_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_blinkt_led_0_avs_s0_writedata;   // mm_interconnect_0:blinkt_led_0_avs_s0_writedata -> blinkt_led_0:avs_s0_writedata
	wire         bytes_to_packets_out_packets_stream_valid;         // bytes_to_packets:out_valid -> avalon_st_adapter:in_0_valid
	wire   [7:0] bytes_to_packets_out_packets_stream_data;          // bytes_to_packets:out_data -> avalon_st_adapter:in_0_data
	wire         bytes_to_packets_out_packets_stream_ready;         // avalon_st_adapter:in_0_ready -> bytes_to_packets:out_ready
	wire   [7:0] bytes_to_packets_out_packets_stream_channel;       // bytes_to_packets:out_channel -> avalon_st_adapter:in_0_channel
	wire         bytes_to_packets_out_packets_stream_startofpacket; // bytes_to_packets:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         bytes_to_packets_out_packets_stream_endofpacket;   // bytes_to_packets:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                     // avalon_st_adapter:out_0_valid -> master:in_valid
	wire   [7:0] avalon_st_adapter_out_0_data;                      // avalon_st_adapter:out_0_data -> master:in_data
	wire         avalon_st_adapter_out_0_ready;                     // master:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;             // avalon_st_adapter:out_0_startofpacket -> master:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;               // avalon_st_adapter:out_0_endofpacket -> master:in_endofpacket
	wire         master_out_stream_valid;                           // master:out_valid -> avalon_st_adapter_001:in_0_valid
	wire   [7:0] master_out_stream_data;                            // master:out_data -> avalon_st_adapter_001:in_0_data
	wire         master_out_stream_ready;                           // avalon_st_adapter_001:in_0_ready -> master:out_ready
	wire         master_out_stream_startofpacket;                   // master:out_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire         master_out_stream_endofpacket;                     // master:out_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire         avalon_st_adapter_001_out_0_valid;                 // avalon_st_adapter_001:out_0_valid -> packets_to_bytes:in_valid
	wire   [7:0] avalon_st_adapter_001_out_0_data;                  // avalon_st_adapter_001:out_0_data -> packets_to_bytes:in_data
	wire         avalon_st_adapter_001_out_0_ready;                 // packets_to_bytes:in_ready -> avalon_st_adapter_001:out_0_ready
	wire   [7:0] avalon_st_adapter_001_out_0_channel;               // avalon_st_adapter_001:out_0_channel -> packets_to_bytes:in_channel
	wire         avalon_st_adapter_001_out_0_startofpacket;         // avalon_st_adapter_001:out_0_startofpacket -> packets_to_bytes:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;           // avalon_st_adapter_001:out_0_endofpacket -> packets_to_bytes:in_endofpacket
	wire         rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, blinkt_led_0:reset_reset, bytes_to_packets:reset_n, master:reset_n, mm_interconnect_0:master_clk_reset_reset_bridge_in_reset_reset, packets_to_bytes:reset_n, simple_led_0:reset_reset]

	apa102_led blinkt_led_0 (
		.avs_s0_address     (mm_interconnect_0_blinkt_led_0_avs_s0_address),     // avs_s0.address
		.avs_s0_read        (mm_interconnect_0_blinkt_led_0_avs_s0_read),        //       .read
		.avs_s0_readdata    (mm_interconnect_0_blinkt_led_0_avs_s0_readdata),    //       .readdata
		.avs_s0_write       (mm_interconnect_0_blinkt_led_0_avs_s0_write),       //       .write
		.avs_s0_writedata   (mm_interconnect_0_blinkt_led_0_avs_s0_writedata),   //       .writedata
		.avs_s0_waitrequest (mm_interconnect_0_blinkt_led_0_avs_s0_waitrequest), //       .waitrequest
		.avs_s0_chipselect  (mm_interconnect_0_blinkt_led_0_avs_s0_chipselect),  //       .chipselect
		.clock_clk          (clk_clk),                                           //  clock.clk
		.reset_reset        (rst_controller_reset_out_reset),                    //  reset.reset
		.sclk               (blinkt_led_serial_serial_clk),                      // serial.serial_clk
		.sdo                (blinkt_led_serial_serial_data)                      //       .serial_data
	);

	altera_avalon_st_bytes_to_packets #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) bytes_to_packets (
		.clk               (clk_clk),                                           //                clk.clk
		.reset_n           (~rst_controller_reset_out_reset),                   //          clk_reset.reset_n
		.out_channel       (bytes_to_packets_out_packets_stream_channel),       // out_packets_stream.channel
		.out_ready         (bytes_to_packets_out_packets_stream_ready),         //                   .ready
		.out_valid         (bytes_to_packets_out_packets_stream_valid),         //                   .valid
		.out_data          (bytes_to_packets_out_packets_stream_data),          //                   .data
		.out_startofpacket (bytes_to_packets_out_packets_stream_startofpacket), //                   .startofpacket
		.out_endofpacket   (bytes_to_packets_out_packets_stream_endofpacket),   //                   .endofpacket
		.in_ready          (bytes_to_packets_in_bytes_stream_ready),            //    in_bytes_stream.ready
		.in_valid          (bytes_to_packets_in_bytes_stream_valid),            //                   .valid
		.in_data           (bytes_to_packets_in_bytes_stream_data)              //                   .data
	);

	altera_avalon_packets_to_master #(
		.FAST_VER    (0),
		.FIFO_DEPTHS (2),
		.FIFO_WIDTHU (1)
	) master (
		.clk               (clk_clk),                               //           clk.clk
		.reset_n           (~rst_controller_reset_out_reset),       //     clk_reset.reset_n
		.out_ready         (master_out_stream_ready),               //    out_stream.ready
		.out_valid         (master_out_stream_valid),               //              .valid
		.out_data          (master_out_stream_data),                //              .data
		.out_startofpacket (master_out_stream_startofpacket),       //              .startofpacket
		.out_endofpacket   (master_out_stream_endofpacket),         //              .endofpacket
		.in_ready          (avalon_st_adapter_out_0_ready),         //     in_stream.ready
		.in_valid          (avalon_st_adapter_out_0_valid),         //              .valid
		.in_data           (avalon_st_adapter_out_0_data),          //              .data
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //              .endofpacket
		.address           (master_avalon_master_address),          // avalon_master.address
		.readdata          (master_avalon_master_readdata),         //              .readdata
		.read              (master_avalon_master_read),             //              .read
		.write             (master_avalon_master_write),            //              .write
		.writedata         (master_avalon_master_writedata),        //              .writedata
		.waitrequest       (master_avalon_master_waitrequest),      //              .waitrequest
		.readdatavalid     (master_avalon_master_readdatavalid),    //              .readdatavalid
		.byteenable        (master_avalon_master_byteenable)        //              .byteenable
	);

	altera_avalon_st_packets_to_bytes #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) packets_to_bytes (
		.clk              (clk_clk),                                   //               clk.clk
		.reset_n          (~rst_controller_reset_out_reset),           //         clk_reset.reset_n
		.in_ready         (avalon_st_adapter_001_out_0_ready),         // in_packets_stream.ready
		.in_valid         (avalon_st_adapter_001_out_0_valid),         //                  .valid
		.in_data          (avalon_st_adapter_001_out_0_data),          //                  .data
		.in_channel       (avalon_st_adapter_001_out_0_channel),       //                  .channel
		.in_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //                  .startofpacket
		.in_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //                  .endofpacket
		.out_ready        (packets_to_bytes_out_bytes_stream_ready),   //  out_bytes_stream.ready
		.out_valid        (packets_to_bytes_out_bytes_stream_valid),   //                  .valid
		.out_data         (packets_to_bytes_out_bytes_stream_data)     //                  .data
	);

	simple_led simple_led_0 (
		.avs_s0_address     (mm_interconnect_0_simple_led_0_avs_s0_address),     //      avs_s0.address
		.avs_s0_read        (mm_interconnect_0_simple_led_0_avs_s0_read),        //            .read
		.avs_s0_readdata    (mm_interconnect_0_simple_led_0_avs_s0_readdata),    //            .readdata
		.avs_s0_write       (mm_interconnect_0_simple_led_0_avs_s0_write),       //            .write
		.avs_s0_writedata   (mm_interconnect_0_simple_led_0_avs_s0_writedata),   //            .writedata
		.avs_s0_waitrequest (mm_interconnect_0_simple_led_0_avs_s0_waitrequest), //            .waitrequest
		.avs_s0_chipselect  (mm_interconnect_0_simple_led_0_avs_s0_chipselect),  //            .chipselect
		.clock_clk          (clk_clk),                                           //       clock.clk
		.reset_reset        (rst_controller_reset_out_reset),                    //       reset.reset
		.out_leds           (simple_leds_leds)                                   // conduit_end.leds
	);

	led_example_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                (clk_clk),                                           //                              clk_0_clk.clk
		.master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // master_clk_reset_reset_bridge_in_reset.reset
		.master_avalon_master_address                 (master_avalon_master_address),                      //                   master_avalon_master.address
		.master_avalon_master_waitrequest             (master_avalon_master_waitrequest),                  //                                       .waitrequest
		.master_avalon_master_byteenable              (master_avalon_master_byteenable),                   //                                       .byteenable
		.master_avalon_master_read                    (master_avalon_master_read),                         //                                       .read
		.master_avalon_master_readdata                (master_avalon_master_readdata),                     //                                       .readdata
		.master_avalon_master_readdatavalid           (master_avalon_master_readdatavalid),                //                                       .readdatavalid
		.master_avalon_master_write                   (master_avalon_master_write),                        //                                       .write
		.master_avalon_master_writedata               (master_avalon_master_writedata),                    //                                       .writedata
		.blinkt_led_0_avs_s0_address                  (mm_interconnect_0_blinkt_led_0_avs_s0_address),     //                    blinkt_led_0_avs_s0.address
		.blinkt_led_0_avs_s0_write                    (mm_interconnect_0_blinkt_led_0_avs_s0_write),       //                                       .write
		.blinkt_led_0_avs_s0_read                     (mm_interconnect_0_blinkt_led_0_avs_s0_read),        //                                       .read
		.blinkt_led_0_avs_s0_readdata                 (mm_interconnect_0_blinkt_led_0_avs_s0_readdata),    //                                       .readdata
		.blinkt_led_0_avs_s0_writedata                (mm_interconnect_0_blinkt_led_0_avs_s0_writedata),   //                                       .writedata
		.blinkt_led_0_avs_s0_waitrequest              (mm_interconnect_0_blinkt_led_0_avs_s0_waitrequest), //                                       .waitrequest
		.blinkt_led_0_avs_s0_chipselect               (mm_interconnect_0_blinkt_led_0_avs_s0_chipselect),  //                                       .chipselect
		.simple_led_0_avs_s0_address                  (mm_interconnect_0_simple_led_0_avs_s0_address),     //                    simple_led_0_avs_s0.address
		.simple_led_0_avs_s0_write                    (mm_interconnect_0_simple_led_0_avs_s0_write),       //                                       .write
		.simple_led_0_avs_s0_read                     (mm_interconnect_0_simple_led_0_avs_s0_read),        //                                       .read
		.simple_led_0_avs_s0_readdata                 (mm_interconnect_0_simple_led_0_avs_s0_readdata),    //                                       .readdata
		.simple_led_0_avs_s0_writedata                (mm_interconnect_0_simple_led_0_avs_s0_writedata),   //                                       .writedata
		.simple_led_0_avs_s0_waitrequest              (mm_interconnect_0_simple_led_0_avs_s0_waitrequest), //                                       .waitrequest
		.simple_led_0_avs_s0_chipselect               (mm_interconnect_0_simple_led_0_avs_s0_chipselect)   //                                       .chipselect
	);

	led_example_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (8),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                    // in_rst_0.reset
		.in_0_data           (bytes_to_packets_out_packets_stream_data),          //     in_0.data
		.in_0_valid          (bytes_to_packets_out_packets_stream_valid),         //         .valid
		.in_0_ready          (bytes_to_packets_out_packets_stream_ready),         //         .ready
		.in_0_startofpacket  (bytes_to_packets_out_packets_stream_startofpacket), //         .startofpacket
		.in_0_endofpacket    (bytes_to_packets_out_packets_stream_endofpacket),   //         .endofpacket
		.in_0_channel        (bytes_to_packets_out_packets_stream_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                      //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                     //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                     //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),             //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                //         .endofpacket
	);

	led_example_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (8),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (master_out_stream_data),                    //     in_0.data
		.in_0_valid          (master_out_stream_valid),                   //         .valid
		.in_0_ready          (master_out_stream_ready),                   //         .ready
		.in_0_startofpacket  (master_out_stream_startofpacket),           //         .startofpacket
		.in_0_endofpacket    (master_out_stream_endofpacket),             //         .endofpacket
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_channel       (avalon_st_adapter_001_out_0_channel)        //         .channel
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
