// avalon_fast_serial.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module avalon_fast_serial (
		input  wire       clk_clk,                //              clk.clk
		output wire       in_bytes_stream_ready,  //  in_bytes_stream.ready
		input  wire       in_bytes_stream_valid,  //                 .valid
		input  wire [7:0] in_bytes_stream_data,   //                 .data
		output wire [7:0] led_gpio_led,           //         led_gpio.led
		input  wire       out_bytes_stream_ready, // out_bytes_stream.ready
		output wire       out_bytes_stream_valid, //                 .valid
		output wire [7:0] out_bytes_stream_data,  //                 .data
		input  wire       reset_reset_n           //            reset.reset_n
	);

	wire  [31:0] master_avalon_master_readdata;                         // mm_interconnect_0:master_avalon_master_readdata -> master:readdata
	wire         master_avalon_master_waitrequest;                      // mm_interconnect_0:master_avalon_master_waitrequest -> master:waitrequest
	wire  [31:0] master_avalon_master_address;                          // master:address -> mm_interconnect_0:master_avalon_master_address
	wire         master_avalon_master_read;                             // master:read -> mm_interconnect_0:master_avalon_master_read
	wire   [3:0] master_avalon_master_byteenable;                       // master:byteenable -> mm_interconnect_0:master_avalon_master_byteenable
	wire         master_avalon_master_readdatavalid;                    // mm_interconnect_0:master_avalon_master_readdatavalid -> master:readdatavalid
	wire         master_avalon_master_write;                            // master:write -> mm_interconnect_0:master_avalon_master_write
	wire  [31:0] master_avalon_master_writedata;                        // master:writedata -> mm_interconnect_0:master_avalon_master_writedata
	wire         riscv_pico_0_avm_m0_chipselect;                        // riscv_pico_0:avm_m0_chipselect -> mm_interconnect_0:riscv_pico_0_avm_m0_chipselect
	wire         riscv_pico_0_avm_m0_waitrequest;                       // mm_interconnect_0:riscv_pico_0_avm_m0_waitrequest -> riscv_pico_0:avm_m0_waitrequest
	wire  [31:0] riscv_pico_0_avm_m0_readdata;                          // mm_interconnect_0:riscv_pico_0_avm_m0_readdata -> riscv_pico_0:avm_m0_readdata
	wire  [15:0] riscv_pico_0_avm_m0_address;                           // riscv_pico_0:avm_m0_address -> mm_interconnect_0:riscv_pico_0_avm_m0_address
	wire         riscv_pico_0_avm_m0_read;                              // riscv_pico_0:avm_m0_read -> mm_interconnect_0:riscv_pico_0_avm_m0_read
	wire         riscv_pico_0_avm_m0_readdatavalid;                     // mm_interconnect_0:riscv_pico_0_avm_m0_readdatavalid -> riscv_pico_0:avm_m0_readdatavalid
	wire         riscv_pico_0_avm_m0_write;                             // riscv_pico_0:avm_m0_write -> mm_interconnect_0:riscv_pico_0_avm_m0_write
	wire  [31:0] riscv_pico_0_avm_m0_writedata;                         // riscv_pico_0:avm_m0_writedata -> mm_interconnect_0:riscv_pico_0_avm_m0_writedata
	wire         mm_interconnect_0_led_gpio_slave_avs_s0_chipselect;    // mm_interconnect_0:led_gpio_slave_avs_s0_chipselect -> led_gpio_slave:avs_s0_chipselect
	wire         mm_interconnect_0_led_gpio_slave_avs_s0_waitrequest;   // led_gpio_slave:avs_s0_waitrequest -> mm_interconnect_0:led_gpio_slave_avs_s0_waitrequest
	wire   [3:0] mm_interconnect_0_led_gpio_slave_avs_s0_address;       // mm_interconnect_0:led_gpio_slave_avs_s0_address -> led_gpio_slave:avs_s0_address
	wire         mm_interconnect_0_led_gpio_slave_avs_s0_write;         // mm_interconnect_0:led_gpio_slave_avs_s0_write -> led_gpio_slave:avs_s0_write
	wire  [31:0] mm_interconnect_0_led_gpio_slave_avs_s0_writedata;     // mm_interconnect_0:led_gpio_slave_avs_s0_writedata -> led_gpio_slave:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata; // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;      // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;        // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire         mm_interconnect_0_onchip_memory2_0_s1_debugaccess;     // mm_interconnect_0:onchip_memory2_0_s1_debugaccess -> onchip_memory2_0:debugaccess
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;         // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;      // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;           // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;       // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;           // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] riscv_pico_0_inr_irq0_irq;                             // irq_mapper:sender_irq -> riscv_pico_0:inr_irq0_irq
	wire         in_bytes_to_packets_out_packets_stream_valid;          // in_bytes_to_packets:out_valid -> avalon_st_adapter:in_0_valid
	wire   [7:0] in_bytes_to_packets_out_packets_stream_data;           // in_bytes_to_packets:out_data -> avalon_st_adapter:in_0_data
	wire         in_bytes_to_packets_out_packets_stream_ready;          // avalon_st_adapter:in_0_ready -> in_bytes_to_packets:out_ready
	wire   [7:0] in_bytes_to_packets_out_packets_stream_channel;        // in_bytes_to_packets:out_channel -> avalon_st_adapter:in_0_channel
	wire         in_bytes_to_packets_out_packets_stream_startofpacket;  // in_bytes_to_packets:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         in_bytes_to_packets_out_packets_stream_endofpacket;    // in_bytes_to_packets:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                         // avalon_st_adapter:out_0_valid -> master:in_valid
	wire   [7:0] avalon_st_adapter_out_0_data;                          // avalon_st_adapter:out_0_data -> master:in_data
	wire         avalon_st_adapter_out_0_ready;                         // master:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                 // avalon_st_adapter:out_0_startofpacket -> master:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                   // avalon_st_adapter:out_0_endofpacket -> master:in_endofpacket
	wire         master_out_stream_valid;                               // master:out_valid -> avalon_st_adapter_001:in_0_valid
	wire   [7:0] master_out_stream_data;                                // master:out_data -> avalon_st_adapter_001:in_0_data
	wire         master_out_stream_ready;                               // avalon_st_adapter_001:in_0_ready -> master:out_ready
	wire         master_out_stream_startofpacket;                       // master:out_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire         master_out_stream_endofpacket;                         // master:out_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire         avalon_st_adapter_001_out_0_valid;                     // avalon_st_adapter_001:out_0_valid -> out_packets_to_bytes:in_valid
	wire   [7:0] avalon_st_adapter_001_out_0_data;                      // avalon_st_adapter_001:out_0_data -> out_packets_to_bytes:in_data
	wire         avalon_st_adapter_001_out_0_ready;                     // out_packets_to_bytes:in_ready -> avalon_st_adapter_001:out_0_ready
	wire   [7:0] avalon_st_adapter_001_out_0_channel;                   // avalon_st_adapter_001:out_0_channel -> out_packets_to_bytes:in_channel
	wire         avalon_st_adapter_001_out_0_startofpacket;             // avalon_st_adapter_001:out_0_startofpacket -> out_packets_to_bytes:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;               // avalon_st_adapter_001:out_0_endofpacket -> out_packets_to_bytes:in_endofpacket
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, in_bytes_to_packets:reset_n, irq_mapper:reset, led_gpio_slave:reset_reset, master:reset_n, mm_interconnect_0:master_clk_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, out_packets_to_bytes:reset_n, riscv_pico_0:reset_reset, rst_translator:in_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	altera_avalon_st_bytes_to_packets #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) in_bytes_to_packets (
		.clk               (clk_clk),                                              //                clk.clk
		.reset_n           (~rst_controller_reset_out_reset),                      //          clk_reset.reset_n
		.out_channel       (in_bytes_to_packets_out_packets_stream_channel),       // out_packets_stream.channel
		.out_ready         (in_bytes_to_packets_out_packets_stream_ready),         //                   .ready
		.out_valid         (in_bytes_to_packets_out_packets_stream_valid),         //                   .valid
		.out_data          (in_bytes_to_packets_out_packets_stream_data),          //                   .data
		.out_startofpacket (in_bytes_to_packets_out_packets_stream_startofpacket), //                   .startofpacket
		.out_endofpacket   (in_bytes_to_packets_out_packets_stream_endofpacket),   //                   .endofpacket
		.in_ready          (in_bytes_stream_ready),                                //    in_bytes_stream.ready
		.in_valid          (in_bytes_stream_valid),                                //                   .valid
		.in_data           (in_bytes_stream_data)                                  //                   .data
	);

	led_gpio led_gpio_slave (
		.avs_s0_address     (mm_interconnect_0_led_gpio_slave_avs_s0_address),     //  avs_s0.address
		.avs_s0_write       (mm_interconnect_0_led_gpio_slave_avs_s0_write),       //        .write
		.avs_s0_writedata   (mm_interconnect_0_led_gpio_slave_avs_s0_writedata),   //        .writedata
		.avs_s0_waitrequest (mm_interconnect_0_led_gpio_slave_avs_s0_waitrequest), //        .waitrequest
		.avs_s0_chipselect  (mm_interconnect_0_led_gpio_slave_avs_s0_chipselect),  //        .chipselect
		.clock_clk          (clk_clk),                                             //   clock.clk
		.reset_reset        (rst_controller_reset_out_reset),                      //   reset.reset
		.LED                (led_gpio_led)                                         // conduit.led
	);

	altera_avalon_packets_to_master #(
		.FAST_VER    (0),
		.FIFO_DEPTHS (2),
		.FIFO_WIDTHU (1)
	) master (
		.clk               (clk_clk),                               //           clk.clk
		.reset_n           (~rst_controller_reset_out_reset),       //     clk_reset.reset_n
		.out_ready         (master_out_stream_ready),               //    out_stream.ready
		.out_valid         (master_out_stream_valid),               //              .valid
		.out_data          (master_out_stream_data),                //              .data
		.out_startofpacket (master_out_stream_startofpacket),       //              .startofpacket
		.out_endofpacket   (master_out_stream_endofpacket),         //              .endofpacket
		.in_ready          (avalon_st_adapter_out_0_ready),         //     in_stream.ready
		.in_valid          (avalon_st_adapter_out_0_valid),         //              .valid
		.in_data           (avalon_st_adapter_out_0_data),          //              .data
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //              .endofpacket
		.address           (master_avalon_master_address),          // avalon_master.address
		.readdata          (master_avalon_master_readdata),         //              .readdata
		.read              (master_avalon_master_read),             //              .read
		.write             (master_avalon_master_write),            //              .write
		.writedata         (master_avalon_master_writedata),        //              .writedata
		.waitrequest       (master_avalon_master_waitrequest),      //              .waitrequest
		.readdatavalid     (master_avalon_master_readdatavalid),    //              .readdatavalid
		.byteenable        (master_avalon_master_byteenable)        //              .byteenable
	);

	avalon_fast_serial_onchip_memory2_0 onchip_memory2_0 (
		.clk         (clk_clk),                                           //   clk1.clk
		.address     (mm_interconnect_0_onchip_memory2_0_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_onchip_memory2_0_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_onchip_memory2_0_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory2_0_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_onchip_memory2_0_s1_write),       //       .write
		.readdata    (mm_interconnect_0_onchip_memory2_0_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory2_0_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory2_0_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),                    // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),                //       .reset_req
		.freeze      (1'b0)                                               // (terminated)
	);

	altera_avalon_st_packets_to_bytes #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) out_packets_to_bytes (
		.clk              (clk_clk),                                   //               clk.clk
		.reset_n          (~rst_controller_reset_out_reset),           //         clk_reset.reset_n
		.in_ready         (avalon_st_adapter_001_out_0_ready),         // in_packets_stream.ready
		.in_valid         (avalon_st_adapter_001_out_0_valid),         //                  .valid
		.in_data          (avalon_st_adapter_001_out_0_data),          //                  .data
		.in_channel       (avalon_st_adapter_001_out_0_channel),       //                  .channel
		.in_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //                  .startofpacket
		.in_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //                  .endofpacket
		.out_ready        (out_bytes_stream_ready),                    //  out_bytes_stream.ready
		.out_valid        (out_bytes_stream_valid),                    //                  .valid
		.out_data         (out_bytes_stream_data)                      //                  .data
	);

	riscv_pico riscv_pico_0 (
		.avm_m0_address       (riscv_pico_0_avm_m0_address),       //   avm_m0.address
		.avm_m0_read          (riscv_pico_0_avm_m0_read),          //         .read
		.avm_m0_waitrequest   (riscv_pico_0_avm_m0_waitrequest),   //         .waitrequest
		.avm_m0_readdata      (riscv_pico_0_avm_m0_readdata),      //         .readdata
		.avm_m0_readdatavalid (riscv_pico_0_avm_m0_readdatavalid), //         .readdatavalid
		.avm_m0_write         (riscv_pico_0_avm_m0_write),         //         .write
		.avm_m0_writedata     (riscv_pico_0_avm_m0_writedata),     //         .writedata
		.avm_m0_chipselect    (riscv_pico_0_avm_m0_chipselect),    //         .chipselect
		.clock_clk            (clk_clk),                           //    clock.clk
		.reset_reset          (rst_controller_reset_out_reset),    //    reset.reset
		.inr_irq0_irq         (riscv_pico_0_inr_irq0_irq)          // inr_irq0.irq
	);

	avalon_fast_serial_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	avalon_fast_serial_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                (clk_clk),                                               //                              clk_0_clk.clk
		.master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // master_clk_reset_reset_bridge_in_reset.reset
		.master_avalon_master_address                 (master_avalon_master_address),                          //                   master_avalon_master.address
		.master_avalon_master_waitrequest             (master_avalon_master_waitrequest),                      //                                       .waitrequest
		.master_avalon_master_byteenable              (master_avalon_master_byteenable),                       //                                       .byteenable
		.master_avalon_master_read                    (master_avalon_master_read),                             //                                       .read
		.master_avalon_master_readdata                (master_avalon_master_readdata),                         //                                       .readdata
		.master_avalon_master_readdatavalid           (master_avalon_master_readdatavalid),                    //                                       .readdatavalid
		.master_avalon_master_write                   (master_avalon_master_write),                            //                                       .write
		.master_avalon_master_writedata               (master_avalon_master_writedata),                        //                                       .writedata
		.riscv_pico_0_avm_m0_address                  (riscv_pico_0_avm_m0_address),                           //                    riscv_pico_0_avm_m0.address
		.riscv_pico_0_avm_m0_waitrequest              (riscv_pico_0_avm_m0_waitrequest),                       //                                       .waitrequest
		.riscv_pico_0_avm_m0_chipselect               (riscv_pico_0_avm_m0_chipselect),                        //                                       .chipselect
		.riscv_pico_0_avm_m0_read                     (riscv_pico_0_avm_m0_read),                              //                                       .read
		.riscv_pico_0_avm_m0_readdata                 (riscv_pico_0_avm_m0_readdata),                          //                                       .readdata
		.riscv_pico_0_avm_m0_readdatavalid            (riscv_pico_0_avm_m0_readdatavalid),                     //                                       .readdatavalid
		.riscv_pico_0_avm_m0_write                    (riscv_pico_0_avm_m0_write),                             //                                       .write
		.riscv_pico_0_avm_m0_writedata                (riscv_pico_0_avm_m0_writedata),                         //                                       .writedata
		.led_gpio_slave_avs_s0_address                (mm_interconnect_0_led_gpio_slave_avs_s0_address),       //                  led_gpio_slave_avs_s0.address
		.led_gpio_slave_avs_s0_write                  (mm_interconnect_0_led_gpio_slave_avs_s0_write),         //                                       .write
		.led_gpio_slave_avs_s0_writedata              (mm_interconnect_0_led_gpio_slave_avs_s0_writedata),     //                                       .writedata
		.led_gpio_slave_avs_s0_waitrequest            (mm_interconnect_0_led_gpio_slave_avs_s0_waitrequest),   //                                       .waitrequest
		.led_gpio_slave_avs_s0_chipselect             (mm_interconnect_0_led_gpio_slave_avs_s0_chipselect),    //                                       .chipselect
		.onchip_memory2_0_s1_address                  (mm_interconnect_0_onchip_memory2_0_s1_address),         //                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                    (mm_interconnect_0_onchip_memory2_0_s1_write),           //                                       .write
		.onchip_memory2_0_s1_readdata                 (mm_interconnect_0_onchip_memory2_0_s1_readdata),        //                                       .readdata
		.onchip_memory2_0_s1_writedata                (mm_interconnect_0_onchip_memory2_0_s1_writedata),       //                                       .writedata
		.onchip_memory2_0_s1_byteenable               (mm_interconnect_0_onchip_memory2_0_s1_byteenable),      //                                       .byteenable
		.onchip_memory2_0_s1_chipselect               (mm_interconnect_0_onchip_memory2_0_s1_chipselect),      //                                       .chipselect
		.onchip_memory2_0_s1_clken                    (mm_interconnect_0_onchip_memory2_0_s1_clken),           //                                       .clken
		.onchip_memory2_0_s1_debugaccess              (mm_interconnect_0_onchip_memory2_0_s1_debugaccess),     //                                       .debugaccess
		.sysid_qsys_0_control_slave_address           (mm_interconnect_0_sysid_qsys_0_control_slave_address),  //             sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata          (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)  //                                       .readdata
	);

	avalon_fast_serial_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (riscv_pico_0_inr_irq0_irq)       //    sender.irq
	);

	avalon_fast_serial_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (8),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                              // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                       // in_rst_0.reset
		.in_0_data           (in_bytes_to_packets_out_packets_stream_data),          //     in_0.data
		.in_0_valid          (in_bytes_to_packets_out_packets_stream_valid),         //         .valid
		.in_0_ready          (in_bytes_to_packets_out_packets_stream_ready),         //         .ready
		.in_0_startofpacket  (in_bytes_to_packets_out_packets_stream_startofpacket), //         .startofpacket
		.in_0_endofpacket    (in_bytes_to_packets_out_packets_stream_endofpacket),   //         .endofpacket
		.in_0_channel        (in_bytes_to_packets_out_packets_stream_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                         //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                        //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                        //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                   //         .endofpacket
	);

	avalon_fast_serial_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (8),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (master_out_stream_data),                    //     in_0.data
		.in_0_valid          (master_out_stream_valid),                   //         .valid
		.in_0_ready          (master_out_stream_ready),                   //         .ready
		.in_0_startofpacket  (master_out_stream_startofpacket),           //         .startofpacket
		.in_0_endofpacket    (master_out_stream_endofpacket),             //         .endofpacket
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_channel       (avalon_st_adapter_001_out_0_channel)        //         .channel
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
